-- Copyright (C) 2021  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- PROGRAM		"Quartus Prime"
-- VERSION		"Version 21.1.0 Build 842 10/21/2021 SJ Lite Edition"
-- CREATED		"Sun Sep 15 18:44:55 2024"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY display IS 
	PORT
	(
		B1 :  IN  STD_LOGIC;
		B2 :  IN  STD_LOGIC;
		B3 :  IN  STD_LOGIC;
		B4 :  IN  STD_LOGIC;
		A :  OUT  STD_LOGIC;
		B :  OUT  STD_LOGIC;
		C :  OUT  STD_LOGIC;
		D :  OUT  STD_LOGIC;
		E :  OUT  STD_LOGIC;
		F :  OUT  STD_LOGIC;
		G :  OUT  STD_LOGIC
	);
END display;

ARCHITECTURE bdf_type OF display IS 

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_35 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_47 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_48 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_49 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_53 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_54 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_55 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_56 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_57 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_58 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_59 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_60 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_61 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_62 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_63 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_64 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_65 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_66 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_67 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_68 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_69 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_70 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_71 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_72 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_73 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_74 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_75 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_76 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_77 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_78 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_79 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_80 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_81 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_82 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_83 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_84 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_85 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_86 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_87 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_88 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_89 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_90 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_91 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_92 :  STD_LOGIC;


BEGIN 



SYNTHESIZED_WIRE_60 <= NOT(B4);



SYNTHESIZED_WIRE_1 <= NOT(B4);



SYNTHESIZED_WIRE_9 <= SYNTHESIZED_WIRE_0 AND SYNTHESIZED_WIRE_1;


G <= NOT(SYNTHESIZED_WIRE_2);



SYNTHESIZED_WIRE_10 <= B1 AND SYNTHESIZED_WIRE_3 AND SYNTHESIZED_WIRE_4;


SYNTHESIZED_WIRE_11 <= SYNTHESIZED_WIRE_5 AND B2 AND B4;


SYNTHESIZED_WIRE_12 <= SYNTHESIZED_WIRE_6 OR SYNTHESIZED_WIRE_7 OR SYNTHESIZED_WIRE_8 OR SYNTHESIZED_WIRE_9 OR SYNTHESIZED_WIRE_10 OR SYNTHESIZED_WIRE_11;


A <= NOT(SYNTHESIZED_WIRE_12);



SYNTHESIZED_WIRE_13 <= NOT(B2);



SYNTHESIZED_WIRE_14 <= NOT(B4);



SYNTHESIZED_WIRE_15 <= NOT(B1);



SYNTHESIZED_WIRE_16 <= NOT(B2);



SYNTHESIZED_WIRE_19 <= NOT(B1);



SYNTHESIZED_WIRE_3 <= NOT(B2);



SYNTHESIZED_WIRE_17 <= NOT(B3);



SYNTHESIZED_WIRE_18 <= NOT(B1);



SYNTHESIZED_WIRE_20 <= NOT(B3);



SYNTHESIZED_WIRE_21 <= NOT(B4);



SYNTHESIZED_WIRE_24 <= SYNTHESIZED_WIRE_13 AND SYNTHESIZED_WIRE_14;


SYNTHESIZED_WIRE_27 <= SYNTHESIZED_WIRE_15 AND SYNTHESIZED_WIRE_16;


SYNTHESIZED_WIRE_25 <= B1 AND SYNTHESIZED_WIRE_17 AND B4;


SYNTHESIZED_WIRE_23 <= SYNTHESIZED_WIRE_18 AND B3 AND B4;


SYNTHESIZED_WIRE_22 <= SYNTHESIZED_WIRE_19 AND SYNTHESIZED_WIRE_20 AND SYNTHESIZED_WIRE_21;


SYNTHESIZED_WIRE_26 <= SYNTHESIZED_WIRE_22 OR SYNTHESIZED_WIRE_23;


SYNTHESIZED_WIRE_5 <= NOT(B1);



SYNTHESIZED_WIRE_28 <= SYNTHESIZED_WIRE_24 OR SYNTHESIZED_WIRE_25 OR SYNTHESIZED_WIRE_26 OR SYNTHESIZED_WIRE_27;


B <= NOT(SYNTHESIZED_WIRE_28);



SYNTHESIZED_WIRE_30 <= NOT(B2);



SYNTHESIZED_WIRE_31 <= NOT(B1);



SYNTHESIZED_WIRE_32 <= NOT(B3);



SYNTHESIZED_WIRE_33 <= NOT(B2);



SYNTHESIZED_WIRE_35 <= NOT(B3);



SYNTHESIZED_WIRE_34 <= NOT(B2);



C <= NOT(SYNTHESIZED_WIRE_29);



SYNTHESIZED_WIRE_38 <= B1 AND SYNTHESIZED_WIRE_30;


SYNTHESIZED_WIRE_0 <= NOT(B2);



SYNTHESIZED_WIRE_41 <= SYNTHESIZED_WIRE_31 AND B2;


SYNTHESIZED_WIRE_39 <= SYNTHESIZED_WIRE_32 AND B4;


SYNTHESIZED_WIRE_37 <= SYNTHESIZED_WIRE_33 AND B4;


SYNTHESIZED_WIRE_36 <= SYNTHESIZED_WIRE_34 AND SYNTHESIZED_WIRE_35;


SYNTHESIZED_WIRE_40 <= SYNTHESIZED_WIRE_36 OR SYNTHESIZED_WIRE_37;


SYNTHESIZED_WIRE_29 <= SYNTHESIZED_WIRE_38 OR SYNTHESIZED_WIRE_39 OR SYNTHESIZED_WIRE_40 OR SYNTHESIZED_WIRE_41;


SYNTHESIZED_WIRE_52 <= B1 AND SYNTHESIZED_WIRE_42 AND B4;


SYNTHESIZED_WIRE_53 <= B2 AND SYNTHESIZED_WIRE_43 AND B4;


SYNTHESIZED_WIRE_54 <= B1 AND B2 AND SYNTHESIZED_WIRE_44;


SYNTHESIZED_WIRE_56 <= SYNTHESIZED_WIRE_45 AND B3 AND B4;


SYNTHESIZED_WIRE_82 <= NOT(B1);



SYNTHESIZED_WIRE_55 <= SYNTHESIZED_WIRE_46 AND B3 AND SYNTHESIZED_WIRE_47;


SYNTHESIZED_WIRE_57 <= SYNTHESIZED_WIRE_48 AND SYNTHESIZED_WIRE_49 AND SYNTHESIZED_WIRE_50;


SYNTHESIZED_WIRE_45 <= NOT(B2);



SYNTHESIZED_WIRE_47 <= NOT(B4);



SYNTHESIZED_WIRE_43 <= NOT(B3);



SYNTHESIZED_WIRE_46 <= NOT(B1);



SYNTHESIZED_WIRE_42 <= NOT(B2);



SYNTHESIZED_WIRE_48 <= NOT(B2);



SYNTHESIZED_WIRE_49 <= NOT(B3);



SYNTHESIZED_WIRE_50 <= NOT(B4);



SYNTHESIZED_WIRE_4 <= NOT(B3);



D <= NOT(SYNTHESIZED_WIRE_51);



SYNTHESIZED_WIRE_44 <= NOT(B4);



SYNTHESIZED_WIRE_51 <= SYNTHESIZED_WIRE_52 OR SYNTHESIZED_WIRE_53 OR SYNTHESIZED_WIRE_54 OR SYNTHESIZED_WIRE_55 OR SYNTHESIZED_WIRE_56 OR SYNTHESIZED_WIRE_57;


SYNTHESIZED_WIRE_62 <= NOT(B4);



SYNTHESIZED_WIRE_59 <= NOT(B4);



SYNTHESIZED_WIRE_61 <= NOT(B2);



E <= NOT(SYNTHESIZED_WIRE_58);



SYNTHESIZED_WIRE_63 <= B1 AND B3;


SYNTHESIZED_WIRE_66 <= B1 AND B2;


SYNTHESIZED_WIRE_64 <= B3 AND SYNTHESIZED_WIRE_59;


SYNTHESIZED_WIRE_6 <= B1 AND SYNTHESIZED_WIRE_60;


SYNTHESIZED_WIRE_65 <= SYNTHESIZED_WIRE_61 AND SYNTHESIZED_WIRE_62;


SYNTHESIZED_WIRE_58 <= SYNTHESIZED_WIRE_63 OR SYNTHESIZED_WIRE_64 OR SYNTHESIZED_WIRE_65 OR SYNTHESIZED_WIRE_66;


SYNTHESIZED_WIRE_76 <= B1 AND SYNTHESIZED_WIRE_67;


SYNTHESIZED_WIRE_79 <= B1 AND B3;


SYNTHESIZED_WIRE_77 <= B2 AND SYNTHESIZED_WIRE_68;


SYNTHESIZED_WIRE_75 <= SYNTHESIZED_WIRE_69 AND SYNTHESIZED_WIRE_70;


SYNTHESIZED_WIRE_74 <= SYNTHESIZED_WIRE_71 AND B2 AND SYNTHESIZED_WIRE_72;


SYNTHESIZED_WIRE_68 <= NOT(B4);



SYNTHESIZED_WIRE_67 <= NOT(B2);



SYNTHESIZED_WIRE_8 <= B2 AND B3;


SYNTHESIZED_WIRE_71 <= NOT(B1);



SYNTHESIZED_WIRE_69 <= NOT(B3);



SYNTHESIZED_WIRE_70 <= NOT(B4);



SYNTHESIZED_WIRE_72 <= NOT(B3);



F <= NOT(SYNTHESIZED_WIRE_73);



SYNTHESIZED_WIRE_78 <= SYNTHESIZED_WIRE_74 OR SYNTHESIZED_WIRE_75;


SYNTHESIZED_WIRE_73 <= SYNTHESIZED_WIRE_76 OR SYNTHESIZED_WIRE_77 OR SYNTHESIZED_WIRE_78 OR SYNTHESIZED_WIRE_79;


SYNTHESIZED_WIRE_87 <= B1 AND SYNTHESIZED_WIRE_80;


SYNTHESIZED_WIRE_89 <= B1 AND B4;


SYNTHESIZED_WIRE_88 <= B3 AND SYNTHESIZED_WIRE_81;


SYNTHESIZED_WIRE_7 <= SYNTHESIZED_WIRE_82 AND B3;


SYNTHESIZED_WIRE_90 <= SYNTHESIZED_WIRE_83 AND B3;


SYNTHESIZED_WIRE_91 <= B2 AND SYNTHESIZED_WIRE_84 AND B4;


SYNTHESIZED_WIRE_92 <= SYNTHESIZED_WIRE_85 AND B2 AND SYNTHESIZED_WIRE_86;


SYNTHESIZED_WIRE_80 <= NOT(B2);



SYNTHESIZED_WIRE_81 <= NOT(B4);



SYNTHESIZED_WIRE_84 <= NOT(B3);



SYNTHESIZED_WIRE_83 <= NOT(B2);



SYNTHESIZED_WIRE_85 <= NOT(B1);



SYNTHESIZED_WIRE_86 <= NOT(B4);



SYNTHESIZED_WIRE_2 <= SYNTHESIZED_WIRE_87 OR SYNTHESIZED_WIRE_88 OR SYNTHESIZED_WIRE_89 OR SYNTHESIZED_WIRE_90 OR SYNTHESIZED_WIRE_91 OR SYNTHESIZED_WIRE_92;


END bdf_type;